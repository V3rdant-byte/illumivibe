// SysForLed.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module SysForLed (
		input  wire        clk_clk,                              //                            clk.clk
		output wire [23:0] color_0_export,                       //                        color_0.export
		output wire [23:0] color_1_export,                       //                        color_1.export
		output wire [23:0] color_10_export,                      //                       color_10.export
		output wire [23:0] color_11_export,                      //                       color_11.export
		output wire [23:0] color_2_export,                       //                        color_2.export
		output wire [23:0] color_3_export,                       //                        color_3.export
		output wire [23:0] color_4_export,                       //                        color_4.export
		output wire [23:0] color_5_export,                       //                        color_5.export
		output wire [23:0] color_6_export,                       //                        color_6.export
		output wire [23:0] color_7_export,                       //                        color_7.export
		output wire [23:0] color_8_export,                       //                        color_8.export
		output wire [23:0] color_9_export,                       //                        color_9.export
		input  wire        reset_reset_n,                        //                          reset.reset_n
		output wire        start_external_connection_export,     //      start_external_connection.export
		input  wire        wifi_uart0_external_connection_rxd,   // wifi_uart0_external_connection.rxd
		output wire        wifi_uart0_external_connection_txd,   //                               .txd
		input  wire        wifi_uart0_external_connection_cts_n, //                               .cts_n
		output wire        wifi_uart0_external_connection_rts_n  //                               .rts_n
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [19:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [19:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_color_0_s1_chipselect;                     // mm_interconnect_0:color_0_s1_chipselect -> color_0:chipselect
	wire  [31:0] mm_interconnect_0_color_0_s1_readdata;                       // color_0:readdata -> mm_interconnect_0:color_0_s1_readdata
	wire   [1:0] mm_interconnect_0_color_0_s1_address;                        // mm_interconnect_0:color_0_s1_address -> color_0:address
	wire         mm_interconnect_0_color_0_s1_write;                          // mm_interconnect_0:color_0_s1_write -> color_0:write_n
	wire  [31:0] mm_interconnect_0_color_0_s1_writedata;                      // mm_interconnect_0:color_0_s1_writedata -> color_0:writedata
	wire         mm_interconnect_0_color_1_s1_chipselect;                     // mm_interconnect_0:color_1_s1_chipselect -> color_1:chipselect
	wire  [31:0] mm_interconnect_0_color_1_s1_readdata;                       // color_1:readdata -> mm_interconnect_0:color_1_s1_readdata
	wire   [1:0] mm_interconnect_0_color_1_s1_address;                        // mm_interconnect_0:color_1_s1_address -> color_1:address
	wire         mm_interconnect_0_color_1_s1_write;                          // mm_interconnect_0:color_1_s1_write -> color_1:write_n
	wire  [31:0] mm_interconnect_0_color_1_s1_writedata;                      // mm_interconnect_0:color_1_s1_writedata -> color_1:writedata
	wire         mm_interconnect_0_color_2_s1_chipselect;                     // mm_interconnect_0:color_2_s1_chipselect -> color_2:chipselect
	wire  [31:0] mm_interconnect_0_color_2_s1_readdata;                       // color_2:readdata -> mm_interconnect_0:color_2_s1_readdata
	wire   [1:0] mm_interconnect_0_color_2_s1_address;                        // mm_interconnect_0:color_2_s1_address -> color_2:address
	wire         mm_interconnect_0_color_2_s1_write;                          // mm_interconnect_0:color_2_s1_write -> color_2:write_n
	wire  [31:0] mm_interconnect_0_color_2_s1_writedata;                      // mm_interconnect_0:color_2_s1_writedata -> color_2:writedata
	wire         mm_interconnect_0_color_3_s1_chipselect;                     // mm_interconnect_0:color_3_s1_chipselect -> color_3:chipselect
	wire  [31:0] mm_interconnect_0_color_3_s1_readdata;                       // color_3:readdata -> mm_interconnect_0:color_3_s1_readdata
	wire   [1:0] mm_interconnect_0_color_3_s1_address;                        // mm_interconnect_0:color_3_s1_address -> color_3:address
	wire         mm_interconnect_0_color_3_s1_write;                          // mm_interconnect_0:color_3_s1_write -> color_3:write_n
	wire  [31:0] mm_interconnect_0_color_3_s1_writedata;                      // mm_interconnect_0:color_3_s1_writedata -> color_3:writedata
	wire         mm_interconnect_0_color_4_s1_chipselect;                     // mm_interconnect_0:color_4_s1_chipselect -> color_4:chipselect
	wire  [31:0] mm_interconnect_0_color_4_s1_readdata;                       // color_4:readdata -> mm_interconnect_0:color_4_s1_readdata
	wire   [1:0] mm_interconnect_0_color_4_s1_address;                        // mm_interconnect_0:color_4_s1_address -> color_4:address
	wire         mm_interconnect_0_color_4_s1_write;                          // mm_interconnect_0:color_4_s1_write -> color_4:write_n
	wire  [31:0] mm_interconnect_0_color_4_s1_writedata;                      // mm_interconnect_0:color_4_s1_writedata -> color_4:writedata
	wire         mm_interconnect_0_color_5_s1_chipselect;                     // mm_interconnect_0:color_5_s1_chipselect -> color_5:chipselect
	wire  [31:0] mm_interconnect_0_color_5_s1_readdata;                       // color_5:readdata -> mm_interconnect_0:color_5_s1_readdata
	wire   [1:0] mm_interconnect_0_color_5_s1_address;                        // mm_interconnect_0:color_5_s1_address -> color_5:address
	wire         mm_interconnect_0_color_5_s1_write;                          // mm_interconnect_0:color_5_s1_write -> color_5:write_n
	wire  [31:0] mm_interconnect_0_color_5_s1_writedata;                      // mm_interconnect_0:color_5_s1_writedata -> color_5:writedata
	wire         mm_interconnect_0_color_6_s1_chipselect;                     // mm_interconnect_0:color_6_s1_chipselect -> color_6:chipselect
	wire  [31:0] mm_interconnect_0_color_6_s1_readdata;                       // color_6:readdata -> mm_interconnect_0:color_6_s1_readdata
	wire   [1:0] mm_interconnect_0_color_6_s1_address;                        // mm_interconnect_0:color_6_s1_address -> color_6:address
	wire         mm_interconnect_0_color_6_s1_write;                          // mm_interconnect_0:color_6_s1_write -> color_6:write_n
	wire  [31:0] mm_interconnect_0_color_6_s1_writedata;                      // mm_interconnect_0:color_6_s1_writedata -> color_6:writedata
	wire         mm_interconnect_0_color_7_s1_chipselect;                     // mm_interconnect_0:color_7_s1_chipselect -> color_7:chipselect
	wire  [31:0] mm_interconnect_0_color_7_s1_readdata;                       // color_7:readdata -> mm_interconnect_0:color_7_s1_readdata
	wire   [1:0] mm_interconnect_0_color_7_s1_address;                        // mm_interconnect_0:color_7_s1_address -> color_7:address
	wire         mm_interconnect_0_color_7_s1_write;                          // mm_interconnect_0:color_7_s1_write -> color_7:write_n
	wire  [31:0] mm_interconnect_0_color_7_s1_writedata;                      // mm_interconnect_0:color_7_s1_writedata -> color_7:writedata
	wire         mm_interconnect_0_color_8_s1_chipselect;                     // mm_interconnect_0:color_8_s1_chipselect -> color_8:chipselect
	wire  [31:0] mm_interconnect_0_color_8_s1_readdata;                       // color_8:readdata -> mm_interconnect_0:color_8_s1_readdata
	wire   [1:0] mm_interconnect_0_color_8_s1_address;                        // mm_interconnect_0:color_8_s1_address -> color_8:address
	wire         mm_interconnect_0_color_8_s1_write;                          // mm_interconnect_0:color_8_s1_write -> color_8:write_n
	wire  [31:0] mm_interconnect_0_color_8_s1_writedata;                      // mm_interconnect_0:color_8_s1_writedata -> color_8:writedata
	wire         mm_interconnect_0_color_9_s1_chipselect;                     // mm_interconnect_0:color_9_s1_chipselect -> color_9:chipselect
	wire  [31:0] mm_interconnect_0_color_9_s1_readdata;                       // color_9:readdata -> mm_interconnect_0:color_9_s1_readdata
	wire   [1:0] mm_interconnect_0_color_9_s1_address;                        // mm_interconnect_0:color_9_s1_address -> color_9:address
	wire         mm_interconnect_0_color_9_s1_write;                          // mm_interconnect_0:color_9_s1_write -> color_9:write_n
	wire  [31:0] mm_interconnect_0_color_9_s1_writedata;                      // mm_interconnect_0:color_9_s1_writedata -> color_9:writedata
	wire         mm_interconnect_0_color_10_s1_chipselect;                    // mm_interconnect_0:color_10_s1_chipselect -> color_10:chipselect
	wire  [31:0] mm_interconnect_0_color_10_s1_readdata;                      // color_10:readdata -> mm_interconnect_0:color_10_s1_readdata
	wire   [1:0] mm_interconnect_0_color_10_s1_address;                       // mm_interconnect_0:color_10_s1_address -> color_10:address
	wire         mm_interconnect_0_color_10_s1_write;                         // mm_interconnect_0:color_10_s1_write -> color_10:write_n
	wire  [31:0] mm_interconnect_0_color_10_s1_writedata;                     // mm_interconnect_0:color_10_s1_writedata -> color_10:writedata
	wire         mm_interconnect_0_color_11_s1_chipselect;                    // mm_interconnect_0:color_11_s1_chipselect -> color_11:chipselect
	wire  [31:0] mm_interconnect_0_color_11_s1_readdata;                      // color_11:readdata -> mm_interconnect_0:color_11_s1_readdata
	wire   [1:0] mm_interconnect_0_color_11_s1_address;                       // mm_interconnect_0:color_11_s1_address -> color_11:address
	wire         mm_interconnect_0_color_11_s1_write;                         // mm_interconnect_0:color_11_s1_write -> color_11:write_n
	wire  [31:0] mm_interconnect_0_color_11_s1_writedata;                     // mm_interconnect_0:color_11_s1_writedata -> color_11:writedata
	wire         mm_interconnect_0_wifi_uart0_s1_chipselect;                  // mm_interconnect_0:wifi_uart0_s1_chipselect -> wifi_uart0:chipselect
	wire  [15:0] mm_interconnect_0_wifi_uart0_s1_readdata;                    // wifi_uart0:readdata -> mm_interconnect_0:wifi_uart0_s1_readdata
	wire   [2:0] mm_interconnect_0_wifi_uart0_s1_address;                     // mm_interconnect_0:wifi_uart0_s1_address -> wifi_uart0:address
	wire         mm_interconnect_0_wifi_uart0_s1_read;                        // mm_interconnect_0:wifi_uart0_s1_read -> wifi_uart0:read_n
	wire         mm_interconnect_0_wifi_uart0_s1_begintransfer;               // mm_interconnect_0:wifi_uart0_s1_begintransfer -> wifi_uart0:begintransfer
	wire         mm_interconnect_0_wifi_uart0_s1_write;                       // mm_interconnect_0:wifi_uart0_s1_write -> wifi_uart0:write_n
	wire  [15:0] mm_interconnect_0_wifi_uart0_s1_writedata;                   // mm_interconnect_0:wifi_uart0_s1_writedata -> wifi_uart0:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_start_s1_chipselect;                       // mm_interconnect_0:start_s1_chipselect -> start:chipselect
	wire  [31:0] mm_interconnect_0_start_s1_readdata;                         // start:readdata -> mm_interconnect_0:start_s1_readdata
	wire   [1:0] mm_interconnect_0_start_s1_address;                          // mm_interconnect_0:start_s1_address -> start:address
	wire         mm_interconnect_0_start_s1_write;                            // mm_interconnect_0:start_s1_write -> start:write_n
	wire  [31:0] mm_interconnect_0_start_s1_writedata;                        // mm_interconnect_0:start_s1_writedata -> start:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                     // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                        // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                          // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                      // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // wifi_uart0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // timer_1:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [color_0:reset_n, color_10:reset_n, color_11:reset_n, color_1:reset_n, color_2:reset_n, color_3:reset_n, color_4:reset_n, color_5:reset_n, color_6:reset_n, color_7:reset_n, color_8:reset_n, color_9:reset_n, jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, start:reset_n, timer_0:reset_n, timer_1:reset_n, wifi_uart0:reset_n]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1

	SysForLed_color_0 color_0 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_0_s1_readdata),   //                    .readdata
		.out_port   (color_0_export)                           // external_connection.export
	);

	SysForLed_color_0 color_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_1_s1_readdata),   //                    .readdata
		.out_port   (color_1_export)                           // external_connection.export
	);

	SysForLed_color_0 color_10 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_color_10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_10_s1_readdata),   //                    .readdata
		.out_port   (color_10_export)                           // external_connection.export
	);

	SysForLed_color_0 color_11 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_color_11_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_11_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_11_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_11_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_11_s1_readdata),   //                    .readdata
		.out_port   (color_11_export)                           // external_connection.export
	);

	SysForLed_color_0 color_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_2_s1_readdata),   //                    .readdata
		.out_port   (color_2_export)                           // external_connection.export
	);

	SysForLed_color_0 color_3 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_3_s1_readdata),   //                    .readdata
		.out_port   (color_3_export)                           // external_connection.export
	);

	SysForLed_color_0 color_4 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_4_s1_readdata),   //                    .readdata
		.out_port   (color_4_export)                           // external_connection.export
	);

	SysForLed_color_0 color_5 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_5_s1_readdata),   //                    .readdata
		.out_port   (color_5_export)                           // external_connection.export
	);

	SysForLed_color_0 color_6 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_6_s1_readdata),   //                    .readdata
		.out_port   (color_6_export)                           // external_connection.export
	);

	SysForLed_color_0 color_7 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_7_s1_readdata),   //                    .readdata
		.out_port   (color_7_export)                           // external_connection.export
	);

	SysForLed_color_0 color_8 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_8_s1_readdata),   //                    .readdata
		.out_port   (color_8_export)                           // external_connection.export
	);

	SysForLed_color_0 color_9 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_color_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_color_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_color_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_color_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_color_9_s1_readdata),   //                    .readdata
		.out_port   (color_9_export)                           // external_connection.export
	);

	SysForLed_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	SysForLed_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	SysForLed_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	SysForLed_start start (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_start_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_s1_readdata),   //                    .readdata
		.out_port   (start_external_connection_export)       // external_connection.export
	);

	SysForLed_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	SysForLed_timer_0 timer_1 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	SysForLed_wifi_uart0 wifi_uart0 (
		.clk           (clk_clk),                                       //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address       (mm_interconnect_0_wifi_uart0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_wifi_uart0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_wifi_uart0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_wifi_uart0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_wifi_uart0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_wifi_uart0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_wifi_uart0_s1_readdata),      //                    .readdata
		.rxd           (wifi_uart0_external_connection_rxd),            // external_connection.export
		.txd           (wifi_uart0_external_connection_txd),            //                    .export
		.cts_n         (wifi_uart0_external_connection_cts_n),          //                    .export
		.rts_n         (wifi_uart0_external_connection_rts_n),          //                    .export
		.irq           (irq_mapper_receiver1_irq)                       //                 irq.irq
	);

	SysForLed_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                              //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                      //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),               //                                         .readdatavalid
		.color_0_s1_address                             (mm_interconnect_0_color_0_s1_address),                        //                               color_0_s1.address
		.color_0_s1_write                               (mm_interconnect_0_color_0_s1_write),                          //                                         .write
		.color_0_s1_readdata                            (mm_interconnect_0_color_0_s1_readdata),                       //                                         .readdata
		.color_0_s1_writedata                           (mm_interconnect_0_color_0_s1_writedata),                      //                                         .writedata
		.color_0_s1_chipselect                          (mm_interconnect_0_color_0_s1_chipselect),                     //                                         .chipselect
		.color_1_s1_address                             (mm_interconnect_0_color_1_s1_address),                        //                               color_1_s1.address
		.color_1_s1_write                               (mm_interconnect_0_color_1_s1_write),                          //                                         .write
		.color_1_s1_readdata                            (mm_interconnect_0_color_1_s1_readdata),                       //                                         .readdata
		.color_1_s1_writedata                           (mm_interconnect_0_color_1_s1_writedata),                      //                                         .writedata
		.color_1_s1_chipselect                          (mm_interconnect_0_color_1_s1_chipselect),                     //                                         .chipselect
		.color_10_s1_address                            (mm_interconnect_0_color_10_s1_address),                       //                              color_10_s1.address
		.color_10_s1_write                              (mm_interconnect_0_color_10_s1_write),                         //                                         .write
		.color_10_s1_readdata                           (mm_interconnect_0_color_10_s1_readdata),                      //                                         .readdata
		.color_10_s1_writedata                          (mm_interconnect_0_color_10_s1_writedata),                     //                                         .writedata
		.color_10_s1_chipselect                         (mm_interconnect_0_color_10_s1_chipselect),                    //                                         .chipselect
		.color_11_s1_address                            (mm_interconnect_0_color_11_s1_address),                       //                              color_11_s1.address
		.color_11_s1_write                              (mm_interconnect_0_color_11_s1_write),                         //                                         .write
		.color_11_s1_readdata                           (mm_interconnect_0_color_11_s1_readdata),                      //                                         .readdata
		.color_11_s1_writedata                          (mm_interconnect_0_color_11_s1_writedata),                     //                                         .writedata
		.color_11_s1_chipselect                         (mm_interconnect_0_color_11_s1_chipselect),                    //                                         .chipselect
		.color_2_s1_address                             (mm_interconnect_0_color_2_s1_address),                        //                               color_2_s1.address
		.color_2_s1_write                               (mm_interconnect_0_color_2_s1_write),                          //                                         .write
		.color_2_s1_readdata                            (mm_interconnect_0_color_2_s1_readdata),                       //                                         .readdata
		.color_2_s1_writedata                           (mm_interconnect_0_color_2_s1_writedata),                      //                                         .writedata
		.color_2_s1_chipselect                          (mm_interconnect_0_color_2_s1_chipselect),                     //                                         .chipselect
		.color_3_s1_address                             (mm_interconnect_0_color_3_s1_address),                        //                               color_3_s1.address
		.color_3_s1_write                               (mm_interconnect_0_color_3_s1_write),                          //                                         .write
		.color_3_s1_readdata                            (mm_interconnect_0_color_3_s1_readdata),                       //                                         .readdata
		.color_3_s1_writedata                           (mm_interconnect_0_color_3_s1_writedata),                      //                                         .writedata
		.color_3_s1_chipselect                          (mm_interconnect_0_color_3_s1_chipselect),                     //                                         .chipselect
		.color_4_s1_address                             (mm_interconnect_0_color_4_s1_address),                        //                               color_4_s1.address
		.color_4_s1_write                               (mm_interconnect_0_color_4_s1_write),                          //                                         .write
		.color_4_s1_readdata                            (mm_interconnect_0_color_4_s1_readdata),                       //                                         .readdata
		.color_4_s1_writedata                           (mm_interconnect_0_color_4_s1_writedata),                      //                                         .writedata
		.color_4_s1_chipselect                          (mm_interconnect_0_color_4_s1_chipselect),                     //                                         .chipselect
		.color_5_s1_address                             (mm_interconnect_0_color_5_s1_address),                        //                               color_5_s1.address
		.color_5_s1_write                               (mm_interconnect_0_color_5_s1_write),                          //                                         .write
		.color_5_s1_readdata                            (mm_interconnect_0_color_5_s1_readdata),                       //                                         .readdata
		.color_5_s1_writedata                           (mm_interconnect_0_color_5_s1_writedata),                      //                                         .writedata
		.color_5_s1_chipselect                          (mm_interconnect_0_color_5_s1_chipselect),                     //                                         .chipselect
		.color_6_s1_address                             (mm_interconnect_0_color_6_s1_address),                        //                               color_6_s1.address
		.color_6_s1_write                               (mm_interconnect_0_color_6_s1_write),                          //                                         .write
		.color_6_s1_readdata                            (mm_interconnect_0_color_6_s1_readdata),                       //                                         .readdata
		.color_6_s1_writedata                           (mm_interconnect_0_color_6_s1_writedata),                      //                                         .writedata
		.color_6_s1_chipselect                          (mm_interconnect_0_color_6_s1_chipselect),                     //                                         .chipselect
		.color_7_s1_address                             (mm_interconnect_0_color_7_s1_address),                        //                               color_7_s1.address
		.color_7_s1_write                               (mm_interconnect_0_color_7_s1_write),                          //                                         .write
		.color_7_s1_readdata                            (mm_interconnect_0_color_7_s1_readdata),                       //                                         .readdata
		.color_7_s1_writedata                           (mm_interconnect_0_color_7_s1_writedata),                      //                                         .writedata
		.color_7_s1_chipselect                          (mm_interconnect_0_color_7_s1_chipselect),                     //                                         .chipselect
		.color_8_s1_address                             (mm_interconnect_0_color_8_s1_address),                        //                               color_8_s1.address
		.color_8_s1_write                               (mm_interconnect_0_color_8_s1_write),                          //                                         .write
		.color_8_s1_readdata                            (mm_interconnect_0_color_8_s1_readdata),                       //                                         .readdata
		.color_8_s1_writedata                           (mm_interconnect_0_color_8_s1_writedata),                      //                                         .writedata
		.color_8_s1_chipselect                          (mm_interconnect_0_color_8_s1_chipselect),                     //                                         .chipselect
		.color_9_s1_address                             (mm_interconnect_0_color_9_s1_address),                        //                               color_9_s1.address
		.color_9_s1_write                               (mm_interconnect_0_color_9_s1_write),                          //                                         .write
		.color_9_s1_readdata                            (mm_interconnect_0_color_9_s1_readdata),                       //                                         .readdata
		.color_9_s1_writedata                           (mm_interconnect_0_color_9_s1_writedata),                      //                                         .writedata
		.color_9_s1_chipselect                          (mm_interconnect_0_color_9_s1_chipselect),                     //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.start_s1_address                               (mm_interconnect_0_start_s1_address),                          //                                 start_s1.address
		.start_s1_write                                 (mm_interconnect_0_start_s1_write),                            //                                         .write
		.start_s1_readdata                              (mm_interconnect_0_start_s1_readdata),                         //                                         .readdata
		.start_s1_writedata                             (mm_interconnect_0_start_s1_writedata),                        //                                         .writedata
		.start_s1_chipselect                            (mm_interconnect_0_start_s1_chipselect),                       //                                         .chipselect
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect),                     //                                         .chipselect
		.timer_1_s1_address                             (mm_interconnect_0_timer_1_s1_address),                        //                               timer_1_s1.address
		.timer_1_s1_write                               (mm_interconnect_0_timer_1_s1_write),                          //                                         .write
		.timer_1_s1_readdata                            (mm_interconnect_0_timer_1_s1_readdata),                       //                                         .readdata
		.timer_1_s1_writedata                           (mm_interconnect_0_timer_1_s1_writedata),                      //                                         .writedata
		.timer_1_s1_chipselect                          (mm_interconnect_0_timer_1_s1_chipselect),                     //                                         .chipselect
		.wifi_uart0_s1_address                          (mm_interconnect_0_wifi_uart0_s1_address),                     //                            wifi_uart0_s1.address
		.wifi_uart0_s1_write                            (mm_interconnect_0_wifi_uart0_s1_write),                       //                                         .write
		.wifi_uart0_s1_read                             (mm_interconnect_0_wifi_uart0_s1_read),                        //                                         .read
		.wifi_uart0_s1_readdata                         (mm_interconnect_0_wifi_uart0_s1_readdata),                    //                                         .readdata
		.wifi_uart0_s1_writedata                        (mm_interconnect_0_wifi_uart0_s1_writedata),                   //                                         .writedata
		.wifi_uart0_s1_begintransfer                    (mm_interconnect_0_wifi_uart0_s1_begintransfer),               //                                         .begintransfer
		.wifi_uart0_s1_chipselect                       (mm_interconnect_0_wifi_uart0_s1_chipselect)                   //                                         .chipselect
	);

	SysForLed_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
